/*

Copyright (c) 2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`timescale 1ns / 1ps

/*
 * AXI4 width adapter
 */
module axi_adapter #(
   // Width of address bus in bits
   parameter ADDR_WIDTH           = 32,
   // Width of input (slave) interface data bus in bits
   parameter S_DATA_WIDTH         = 32,
   // Width of input (slave) interface wstrb (width of data bus in words)
   parameter S_STRB_WIDTH         = (S_DATA_WIDTH / 8),
   // Width of output (master) interface data bus in bits
   parameter M_DATA_WIDTH         = 32,
   // Width of output (master) interface wstrb (width of data bus in words)
   parameter M_STRB_WIDTH         = (M_DATA_WIDTH / 8),
   // Width of ID signal
   parameter ID_WIDTH             = 8,
   // Propagate awuser signal
   parameter AWUSER_ENABLE        = 0,
   // Width of awuser signal
   parameter AWUSER_WIDTH         = 1,
   // Propagate wuser signal
   parameter WUSER_ENABLE         = 0,
   // Width of wuser signal
   parameter WUSER_WIDTH          = 1,
   // Propagate buser signal
   parameter BUSER_ENABLE         = 0,
   // Width of buser signal
   parameter BUSER_WIDTH          = 1,
   // Propagate aruser signal
   parameter ARUSER_ENABLE        = 0,
   // Width of aruser signal
   parameter ARUSER_WIDTH         = 1,
   // Propagate ruser signal
   parameter RUSER_ENABLE         = 0,
   // Width of ruser signal
   parameter RUSER_WIDTH          = 1,
   // When adapting to a wider bus, re-pack full-width burst instead of passing through narrow burst if possible
   parameter CONVERT_BURST        = 1,
   // When adapting to a wider bus, re-pack all bursts instead of passing through narrow burst if possible
   parameter CONVERT_NARROW_BURST = 0,
   // Forward ID through adapter
   parameter FORWARD_ID           = 0
) (
   input wire clk,
   input wire rst,

   /*
     * AXI slave interface
     */
   input  wire [    ID_WIDTH-1:0] s_axi_awid,
   input  wire [  ADDR_WIDTH-1:0] s_axi_awaddr,
   input  wire [             7:0] s_axi_awlen,
   input  wire [             2:0] s_axi_awsize,
   input  wire [             1:0] s_axi_awburst,
   input  wire                    s_axi_awlock,
   input  wire [             3:0] s_axi_awcache,
   input  wire [             2:0] s_axi_awprot,
   input  wire [             3:0] s_axi_awqos,
   input  wire [             3:0] s_axi_awregion,
   input  wire [AWUSER_WIDTH-1:0] s_axi_awuser,
   input  wire                    s_axi_awvalid,
   output wire                    s_axi_awready,
   input  wire [S_DATA_WIDTH-1:0] s_axi_wdata,
   input  wire [S_STRB_WIDTH-1:0] s_axi_wstrb,
   input  wire                    s_axi_wlast,
   input  wire [ WUSER_WIDTH-1:0] s_axi_wuser,
   input  wire                    s_axi_wvalid,
   output wire                    s_axi_wready,
   output wire [    ID_WIDTH-1:0] s_axi_bid,
   output wire [             1:0] s_axi_bresp,
   output wire [ BUSER_WIDTH-1:0] s_axi_buser,
   output wire                    s_axi_bvalid,
   input  wire                    s_axi_bready,
   input  wire [    ID_WIDTH-1:0] s_axi_arid,
   input  wire [  ADDR_WIDTH-1:0] s_axi_araddr,
   input  wire [             7:0] s_axi_arlen,
   input  wire [             2:0] s_axi_arsize,
   input  wire [             1:0] s_axi_arburst,
   input  wire                    s_axi_arlock,
   input  wire [             3:0] s_axi_arcache,
   input  wire [             2:0] s_axi_arprot,
   input  wire [             3:0] s_axi_arqos,
   input  wire [             3:0] s_axi_arregion,
   input  wire [ARUSER_WIDTH-1:0] s_axi_aruser,
   input  wire                    s_axi_arvalid,
   output wire                    s_axi_arready,
   output wire [    ID_WIDTH-1:0] s_axi_rid,
   output wire [S_DATA_WIDTH-1:0] s_axi_rdata,
   output wire [             1:0] s_axi_rresp,
   output wire                    s_axi_rlast,
   output wire [ RUSER_WIDTH-1:0] s_axi_ruser,
   output wire                    s_axi_rvalid,
   input  wire                    s_axi_rready,

   /*
     * AXI master interface
     */
   output wire [    ID_WIDTH-1:0] m_axi_awid,
   output wire [  ADDR_WIDTH-1:0] m_axi_awaddr,
   output wire [             7:0] m_axi_awlen,
   output wire [             2:0] m_axi_awsize,
   output wire [             1:0] m_axi_awburst,
   output wire                    m_axi_awlock,
   output wire [             3:0] m_axi_awcache,
   output wire [             2:0] m_axi_awprot,
   output wire [             3:0] m_axi_awqos,
   output wire [             3:0] m_axi_awregion,
   output wire [AWUSER_WIDTH-1:0] m_axi_awuser,
   output wire                    m_axi_awvalid,
   input  wire                    m_axi_awready,
   output wire [M_DATA_WIDTH-1:0] m_axi_wdata,
   output wire [M_STRB_WIDTH-1:0] m_axi_wstrb,
   output wire                    m_axi_wlast,
   output wire [ WUSER_WIDTH-1:0] m_axi_wuser,
   output wire                    m_axi_wvalid,
   input  wire                    m_axi_wready,
   input  wire [    ID_WIDTH-1:0] m_axi_bid,
   input  wire [             1:0] m_axi_bresp,
   input  wire [ BUSER_WIDTH-1:0] m_axi_buser,
   input  wire                    m_axi_bvalid,
   output wire                    m_axi_bready,
   output wire [    ID_WIDTH-1:0] m_axi_arid,
   output wire [  ADDR_WIDTH-1:0] m_axi_araddr,
   output wire [             7:0] m_axi_arlen,
   output wire [             2:0] m_axi_arsize,
   output wire [             1:0] m_axi_arburst,
   output wire                    m_axi_arlock,
   output wire [             3:0] m_axi_arcache,
   output wire [             2:0] m_axi_arprot,
   output wire [             3:0] m_axi_arqos,
   output wire [             3:0] m_axi_arregion,
   output wire [ARUSER_WIDTH-1:0] m_axi_aruser,
   output wire                    m_axi_arvalid,
   input  wire                    m_axi_arready,
   input  wire [    ID_WIDTH-1:0] m_axi_rid,
   input  wire [M_DATA_WIDTH-1:0] m_axi_rdata,
   input  wire [             1:0] m_axi_rresp,
   input  wire                    m_axi_rlast,
   input  wire [ RUSER_WIDTH-1:0] m_axi_ruser,
   input  wire                    m_axi_rvalid,
   output wire                    m_axi_rready
);

   axi_adapter_wr #(
      .ADDR_WIDTH          (ADDR_WIDTH),
      .S_DATA_WIDTH        (S_DATA_WIDTH),
      .S_STRB_WIDTH        (S_STRB_WIDTH),
      .M_DATA_WIDTH        (M_DATA_WIDTH),
      .M_STRB_WIDTH        (M_STRB_WIDTH),
      .ID_WIDTH            (ID_WIDTH),
      .AWUSER_ENABLE       (AWUSER_ENABLE),
      .AWUSER_WIDTH        (AWUSER_WIDTH),
      .WUSER_ENABLE        (WUSER_ENABLE),
      .WUSER_WIDTH         (WUSER_WIDTH),
      .BUSER_ENABLE        (BUSER_ENABLE),
      .BUSER_WIDTH         (BUSER_WIDTH),
      .CONVERT_BURST       (CONVERT_BURST),
      .CONVERT_NARROW_BURST(CONVERT_NARROW_BURST),
      .FORWARD_ID          (FORWARD_ID)
   ) axi_adapter_wr_inst (
      .clk(clk),
      .rst(rst),

      /*
     * AXI slave interface
     */
      .s_axi_awid    (s_axi_awid),
      .s_axi_awaddr  (s_axi_awaddr),
      .s_axi_awlen   (s_axi_awlen),
      .s_axi_awsize  (s_axi_awsize),
      .s_axi_awburst (s_axi_awburst),
      .s_axi_awlock  (s_axi_awlock),
      .s_axi_awcache (s_axi_awcache),
      .s_axi_awprot  (s_axi_awprot),
      .s_axi_awqos   (s_axi_awqos),
      .s_axi_awregion(s_axi_awregion),
      .s_axi_awuser  (s_axi_awuser),
      .s_axi_awvalid (s_axi_awvalid),
      .s_axi_awready (s_axi_awready),
      .s_axi_wdata   (s_axi_wdata),
      .s_axi_wstrb   (s_axi_wstrb),
      .s_axi_wlast   (s_axi_wlast),
      .s_axi_wuser   (s_axi_wuser),
      .s_axi_wvalid  (s_axi_wvalid),
      .s_axi_wready  (s_axi_wready),
      .s_axi_bid     (s_axi_bid),
      .s_axi_bresp   (s_axi_bresp),
      .s_axi_buser   (s_axi_buser),
      .s_axi_bvalid  (s_axi_bvalid),
      .s_axi_bready  (s_axi_bready),

      /*
     * AXI master interface
     */
      .m_axi_awid    (m_axi_awid),
      .m_axi_awaddr  (m_axi_awaddr),
      .m_axi_awlen   (m_axi_awlen),
      .m_axi_awsize  (m_axi_awsize),
      .m_axi_awburst (m_axi_awburst),
      .m_axi_awlock  (m_axi_awlock),
      .m_axi_awcache (m_axi_awcache),
      .m_axi_awprot  (m_axi_awprot),
      .m_axi_awqos   (m_axi_awqos),
      .m_axi_awregion(m_axi_awregion),
      .m_axi_awuser  (m_axi_awuser),
      .m_axi_awvalid (m_axi_awvalid),
      .m_axi_awready (m_axi_awready),
      .m_axi_wdata   (m_axi_wdata),
      .m_axi_wstrb   (m_axi_wstrb),
      .m_axi_wlast   (m_axi_wlast),
      .m_axi_wuser   (m_axi_wuser),
      .m_axi_wvalid  (m_axi_wvalid),
      .m_axi_wready  (m_axi_wready),
      .m_axi_bid     (m_axi_bid),
      .m_axi_bresp   (m_axi_bresp),
      .m_axi_buser   (m_axi_buser),
      .m_axi_bvalid  (m_axi_bvalid),
      .m_axi_bready  (m_axi_bready)
   );

   axi_adapter_rd #(
      .ADDR_WIDTH          (ADDR_WIDTH),
      .S_DATA_WIDTH        (S_DATA_WIDTH),
      .S_STRB_WIDTH        (S_STRB_WIDTH),
      .M_DATA_WIDTH        (M_DATA_WIDTH),
      .M_STRB_WIDTH        (M_STRB_WIDTH),
      .ID_WIDTH            (ID_WIDTH),
      .ARUSER_ENABLE       (ARUSER_ENABLE),
      .ARUSER_WIDTH        (ARUSER_WIDTH),
      .RUSER_ENABLE        (RUSER_ENABLE),
      .RUSER_WIDTH         (RUSER_WIDTH),
      .CONVERT_BURST       (CONVERT_BURST),
      .CONVERT_NARROW_BURST(CONVERT_NARROW_BURST),
      .FORWARD_ID          (FORWARD_ID)
   ) axi_adapter_rd_inst (
      .clk(clk),
      .rst(rst),

      /*
     * AXI slave interface
     */
      .s_axi_arid    (s_axi_arid),
      .s_axi_araddr  (s_axi_araddr),
      .s_axi_arlen   (s_axi_arlen),
      .s_axi_arsize  (s_axi_arsize),
      .s_axi_arburst (s_axi_arburst),
      .s_axi_arlock  (s_axi_arlock),
      .s_axi_arcache (s_axi_arcache),
      .s_axi_arprot  (s_axi_arprot),
      .s_axi_arqos   (s_axi_arqos),
      .s_axi_arregion(s_axi_arregion),
      .s_axi_aruser  (s_axi_aruser),
      .s_axi_arvalid (s_axi_arvalid),
      .s_axi_arready (s_axi_arready),
      .s_axi_rid     (s_axi_rid),
      .s_axi_rdata   (s_axi_rdata),
      .s_axi_rresp   (s_axi_rresp),
      .s_axi_rlast   (s_axi_rlast),
      .s_axi_ruser   (s_axi_ruser),
      .s_axi_rvalid  (s_axi_rvalid),
      .s_axi_rready  (s_axi_rready),

      /*
     * AXI master interface
     */
      .m_axi_arid    (m_axi_arid),
      .m_axi_araddr  (m_axi_araddr),
      .m_axi_arlen   (m_axi_arlen),
      .m_axi_arsize  (m_axi_arsize),
      .m_axi_arburst (m_axi_arburst),
      .m_axi_arlock  (m_axi_arlock),
      .m_axi_arcache (m_axi_arcache),
      .m_axi_arprot  (m_axi_arprot),
      .m_axi_arqos   (m_axi_arqos),
      .m_axi_arregion(m_axi_arregion),
      .m_axi_aruser  (m_axi_aruser),
      .m_axi_arvalid (m_axi_arvalid),
      .m_axi_arready (m_axi_arready),
      .m_axi_rid     (m_axi_rid),
      .m_axi_rdata   (m_axi_rdata),
      .m_axi_rresp   (m_axi_rresp),
      .m_axi_rlast   (m_axi_rlast),
      .m_axi_ruser   (m_axi_ruser),
      .m_axi_rvalid  (m_axi_rvalid),
      .m_axi_rready  (m_axi_rready)
   );

endmodule
