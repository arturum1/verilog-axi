/*

Copyright (c) 2019 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`timescale 1ns / 1ps

/*
 * AXI4 lite clock domain crossing module
 */
module axil_cdc #(
   // Width of data bus in bits
   parameter DATA_WIDTH = 32,
   // Width of address bus in bits
   parameter ADDR_WIDTH = 32,
   // Width of wstrb (width of data bus in words)
   parameter STRB_WIDTH = (DATA_WIDTH / 8)
) (
   /*
     * AXI lite slave interface
     */
   input  wire                  s_clk,
   input  wire                  s_rst,
   input  wire [ADDR_WIDTH-1:0] s_axil_awaddr,
   input  wire [           2:0] s_axil_awprot,
   input  wire                  s_axil_awvalid,
   output wire                  s_axil_awready,
   input  wire [DATA_WIDTH-1:0] s_axil_wdata,
   input  wire [STRB_WIDTH-1:0] s_axil_wstrb,
   input  wire                  s_axil_wvalid,
   output wire                  s_axil_wready,
   output wire [           1:0] s_axil_bresp,
   output wire                  s_axil_bvalid,
   input  wire                  s_axil_bready,
   input  wire [ADDR_WIDTH-1:0] s_axil_araddr,
   input  wire [           2:0] s_axil_arprot,
   input  wire                  s_axil_arvalid,
   output wire                  s_axil_arready,
   output wire [DATA_WIDTH-1:0] s_axil_rdata,
   output wire [           1:0] s_axil_rresp,
   output wire                  s_axil_rvalid,
   input  wire                  s_axil_rready,

   /*
     * AXI lite master interface
     */
   input  wire                  m_clk,
   input  wire                  m_rst,
   output wire [ADDR_WIDTH-1:0] m_axil_awaddr,
   output wire [           2:0] m_axil_awprot,
   output wire                  m_axil_awvalid,
   input  wire                  m_axil_awready,
   output wire [DATA_WIDTH-1:0] m_axil_wdata,
   output wire [STRB_WIDTH-1:0] m_axil_wstrb,
   output wire                  m_axil_wvalid,
   input  wire                  m_axil_wready,
   input  wire [           1:0] m_axil_bresp,
   input  wire                  m_axil_bvalid,
   output wire                  m_axil_bready,
   output wire [ADDR_WIDTH-1:0] m_axil_araddr,
   output wire [           2:0] m_axil_arprot,
   output wire                  m_axil_arvalid,
   input  wire                  m_axil_arready,
   input  wire [DATA_WIDTH-1:0] m_axil_rdata,
   input  wire [           1:0] m_axil_rresp,
   input  wire                  m_axil_rvalid,
   output wire                  m_axil_rready
);

   axil_cdc_wr #(
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(ADDR_WIDTH),
      .STRB_WIDTH(STRB_WIDTH)
   ) axil_cdc_wr_inst (
      /*
     * AXI lite slave interface
     */
      .s_clk         (s_clk),
      .s_rst         (s_rst),
      .s_axil_awaddr (s_axil_awaddr),
      .s_axil_awprot (s_axil_awprot),
      .s_axil_awvalid(s_axil_awvalid),
      .s_axil_awready(s_axil_awready),
      .s_axil_wdata  (s_axil_wdata),
      .s_axil_wstrb  (s_axil_wstrb),
      .s_axil_wvalid (s_axil_wvalid),
      .s_axil_wready (s_axil_wready),
      .s_axil_bresp  (s_axil_bresp),
      .s_axil_bvalid (s_axil_bvalid),
      .s_axil_bready (s_axil_bready),

      /*
     * AXI lite master interface
     */
      .m_clk         (m_clk),
      .m_rst         (m_rst),
      .m_axil_awaddr (m_axil_awaddr),
      .m_axil_awprot (m_axil_awprot),
      .m_axil_awvalid(m_axil_awvalid),
      .m_axil_awready(m_axil_awready),
      .m_axil_wdata  (m_axil_wdata),
      .m_axil_wstrb  (m_axil_wstrb),
      .m_axil_wvalid (m_axil_wvalid),
      .m_axil_wready (m_axil_wready),
      .m_axil_bresp  (m_axil_bresp),
      .m_axil_bvalid (m_axil_bvalid),
      .m_axil_bready (m_axil_bready)
   );

   axil_cdc_rd #(
      .DATA_WIDTH(DATA_WIDTH),
      .ADDR_WIDTH(ADDR_WIDTH),
      .STRB_WIDTH(STRB_WIDTH)
   ) axil_cdc_rd_inst (
      /*
     * AXI lite slave interface
     */
      .s_clk         (s_clk),
      .s_rst         (s_rst),
      .s_axil_araddr (s_axil_araddr),
      .s_axil_arprot (s_axil_arprot),
      .s_axil_arvalid(s_axil_arvalid),
      .s_axil_arready(s_axil_arready),
      .s_axil_rdata  (s_axil_rdata),
      .s_axil_rresp  (s_axil_rresp),
      .s_axil_rvalid (s_axil_rvalid),
      .s_axil_rready (s_axil_rready),

      /*
     * AXI lite master interface
     */
      .m_clk         (m_clk),
      .m_rst         (m_rst),
      .m_axil_araddr (m_axil_araddr),
      .m_axil_arprot (m_axil_arprot),
      .m_axil_arvalid(m_axil_arvalid),
      .m_axil_arready(m_axil_arready),
      .m_axil_rdata  (m_axil_rdata),
      .m_axil_rresp  (m_axil_rresp),
      .m_axil_rvalid (m_axil_rvalid),
      .m_axil_rready (m_axil_rready)
   );

endmodule
